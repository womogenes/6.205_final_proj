parameter integer INV_SQRT_STAGE_DELAY = 5;
parameter integer INV_SQRT_NR_STAGES = 3;
parameter integer INV_SQRT_DELAY = INV_SQRT_NR_STAGES * INV_SQRT_STAGE_DELAY;
