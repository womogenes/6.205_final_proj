// Normalize a vec3 into a vec3s

module normalize (
  input wire clk,
  input wire rst,

  input vec3 din,
  input wire din_valid,

  output vec3 dout,
  output logic dout_valid
);
  // TODO: normalize module
endmodule
