`default_nettype none

`default_nettype wire
