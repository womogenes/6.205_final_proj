// Convert integers to FP24 and vice versa
// Turn 32-bit integer into FP24

module make_fp24 (
  input wire [31:0] n,
  output fp24 x
);
  
endmodule
