// Addition for 24-bit floating point

module fp24_add (
  input wire clk,
  input wire rst,
  input logic [23:0] a,
  input logic [23:0] b,

  output logic [23:0] sum
);
  // TODO: implement
endmodule
