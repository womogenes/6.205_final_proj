// Vector operations (fp24 vec3 add and multiply)
