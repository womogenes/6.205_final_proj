`default_nettype none

module cpu_top_level (
  input wire clk,
  input wire rst
);

  // Expose some stuff for CPU debugging

endmodule

`default_nettype wire
