`default_nettype none

module object_buffer (
  input wire [7:0] obj_idx,

  output object obj
);
  // Read out objects from memory
  
endmodule

`default_nettype wire
