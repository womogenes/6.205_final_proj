typedef enum logic [2:0] { LW, LH, LHU, LB, LBU, SW, SH, SB } MemFunc;
