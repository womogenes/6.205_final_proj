parameter integer FRAC_WIDTH = 16;
parameter integer FULL_WIDTH = 32;

// ===== NUMBERS + MATH =====
// FIXED-POINT TYPES NOT USED
// typedef logic signed [FULL_WIDTH-1:0] fixed;
// typedef logic signed [FRAC_WIDTH:0] short;     // extra bit for two's complement

typedef struct packed {
  logic sign;
  logic [FP_EXP_BITS-1:0] exp;
  logic [FP_MANT_BITS-1:0] mant;
} fp;

// ===== COLORS =====
typedef struct packed {
  logic [7:0] r;
  logic [7:0] g;
  logic [7:0] b;
} color8;

typedef struct packed {
  fp r;
  fp g;
  fp b;
} fp_color;

// ===== VECTOR TYPES =====
typedef struct packed {
  fp x;
  fp y;
  fp z;
} fp_vec3;

// ===== CAMERA =====
typedef struct packed {
  fp_vec3 origin;
  fp_vec3 forward;
  fp_vec3 right;
  fp_vec3 up;
} camera;

// ===== OBJECTS =====
typedef struct packed {
  fp_color color;           // 72 bits
  fp_color emit_color;      // 72 bits
  fp_color spec_color;      // 72 bits
  fp smoothness;            // 24 bits
  logic [7:0] specular_prob;  // 8 bits
} material;

typedef struct packed {
  logic is_trig;            // 1 bit
  material mat;             // [several] bits
  fp_vec3 [2:0] trig;     // 216 bits
  fp_vec3 trig_norm;      // 72 bits
  fp_vec3 sphere_center;  // 72 bits
  fp sphere_rad_sq;       // 24 bits
  fp sphere_rad_inv;      // 24 bits
} object;
