typedef enum { LW, LH, LHU, LB, LBU, SW, SH, SB } MemFunc;
